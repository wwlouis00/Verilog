module hello_world (
    input a,
    input b,

    output y
);

assign y = a & b;
    
endmodule